module collision_detection (
    input,
    output
);

endmodule