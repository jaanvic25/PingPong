module paddle_movement_tb (
    wire enc1a, enc1b, enc2a, enc2b;
);

endmodule