/* 
August 2024
Jaanvi Chirimar, Josie Chan, Sirrye Pierre

Start the game, reset memory (paddle and ball position, scores)
*/

module init (
    // Player scores
    input wire p1,
    input wire p2,

    // Ball position on LED matrix
    input wire b_x,
    input wire b_y,

    // Paddle 1 position on LED matrix
    input wire p1_x,
    input wire p1_y,

    // Paddle 2 position on LED matrix
    input wire p2_x,
    input wire p2_y
);

endmodule